/////////////////////////////////////////////////////////////////////
// Design unit: 
//            :
// File name  : 
//            :
// Description: control of the interrup
//            :
// Limitations:
//            :
// System     : SystemVerilog IEEE 1800-2005
//            :
// Author     : Letian(Brian) Chen
//
// Revision   : Version 0.0 10/2024
/////////////////////////////////////////////////////////////////////
module interrupt (
    
);
    
endmodule